*** Model Description ***
.param temp=27
.param Wp=0.84
.param Wn=0.36

*** Including sky130 library files ***
.lib "sky130_fd_pr/models/sky130.lib.spice" tt

*** Netlist Description ***
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 w={Wp} l=0.15
XM2 out in 0 0 sky130_fd_pr__nfet_01v8 w={Wn}l=0.15
Cload out 0 50fF
Vdd vdd 0 1.8V
Vin in 0 1.8V

*** Simulation Commands ***
.dc Vin 0 1.8 0.01

.control
let idx=1
let loops=40
let Wp_incr=0.84
let Wn_incr=0.36
let Wp_start=0.84
let Wn_start=0.36*20
set c = " "
let vector_Vm = vector(loops)
let vector_Wp_Wn_ratio = vector(loops)

dowhile idx <= loops
    if (idx <= 20)
        let new_Wn = Wn_start - ((idx-1) * Wn_incr)
        let new_Wp = 0.84
    end
    if (idx >= 21)
        let new_Wn = 0.36
        let new_Wp = Wp_start + ((idx-20) * Wp_incr)
    end

    alterparam Wp=$&new_Wp
    alterparam Wn=$&new_Wn
    reset
    run
    meas dc Vm find V(out) when V(out)=V(in)
    let vector_Vm[idx-1] = Vm
    let vector_Wp_Wn_ratio[idx-1] = ($&new_Wp/ $&new_Wn)
    print ($&new_Wp/ $&new_Wn)
    set c = ( $c dc{$&idx}.V(out) )
    let idx = idx + 1
end

set nolegend
plot $c xlabel 'Vin' ylabel 'Vout'
plot vector_Vm vs vector_Wp_Wn_ratio xlabel 'Wp/Wn' ylabel 'Vm (V)'
*+ xlimit vector_Wp_Wn_ratio[0] vector_Wp_Wn_ratio[39] ylimit vector_Vm[0] vector_Vm[39]
.endc

.end